module And (input a , b , output c );
  c2 cell1 (0,1,0,1,1,1,a ,b,c);
endmodule
