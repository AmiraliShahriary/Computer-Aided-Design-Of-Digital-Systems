module carry_out(input a, b, c ,output o);
    c2 co(0,1,c,1,a,b,a,b,o);
endmodule
