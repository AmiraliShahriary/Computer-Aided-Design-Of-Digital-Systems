module inverter(input a , output b);
  c2 cell1 (1,0,1,0,1,1,a,1,b);

endmodule